-----------------------------------------------------------
-- An LU (logic unit) which is responsible for logical operations in the ALU
-- Author: Aaron Moser
-- Date: 12.01.2019
-----------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity lu is
end entity;

